VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_example
  CLASS BLOCK ;
  FOREIGN tt_um_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 149.980 8.810 158.600 10.610 ;
        RECT 149.980 3.790 151.780 8.810 ;
        RECT 156.800 3.790 158.600 8.810 ;
        RECT 149.980 1.990 158.600 3.790 ;
      LAYER li1 ;
        RECT 150.610 9.650 157.970 9.980 ;
        RECT 150.610 2.950 150.940 9.650 ;
        RECT 152.620 7.640 155.960 7.970 ;
        RECT 152.620 4.960 152.950 7.640 ;
        RECT 153.785 5.795 154.795 6.805 ;
        RECT 155.630 4.960 155.960 7.640 ;
        RECT 152.620 4.630 155.960 4.960 ;
        RECT 157.640 2.950 157.970 9.650 ;
        RECT 150.610 2.620 157.970 2.950 ;
      LAYER mcon ;
        RECT 150.690 9.730 150.860 9.900 ;
        RECT 151.145 9.730 151.315 9.900 ;
        RECT 151.505 9.730 151.675 9.900 ;
        RECT 151.865 9.730 152.035 9.900 ;
        RECT 152.225 9.730 152.395 9.900 ;
        RECT 152.585 9.730 152.755 9.900 ;
        RECT 152.945 9.730 153.115 9.900 ;
        RECT 153.305 9.730 153.475 9.900 ;
        RECT 153.665 9.730 153.835 9.900 ;
        RECT 154.025 9.730 154.195 9.900 ;
        RECT 154.385 9.730 154.555 9.900 ;
        RECT 154.745 9.730 154.915 9.900 ;
        RECT 155.105 9.730 155.275 9.900 ;
        RECT 155.465 9.730 155.635 9.900 ;
        RECT 155.825 9.730 155.995 9.900 ;
        RECT 156.185 9.730 156.355 9.900 ;
        RECT 156.545 9.730 156.715 9.900 ;
        RECT 156.905 9.730 157.075 9.900 ;
        RECT 157.265 9.730 157.435 9.900 ;
        RECT 157.720 9.730 157.890 9.900 ;
        RECT 150.690 9.275 150.860 9.445 ;
        RECT 150.690 8.915 150.860 9.085 ;
        RECT 150.690 8.555 150.860 8.725 ;
        RECT 150.690 8.195 150.860 8.365 ;
        RECT 150.690 7.835 150.860 8.005 ;
        RECT 157.720 9.275 157.890 9.445 ;
        RECT 157.720 8.915 157.890 9.085 ;
        RECT 157.720 8.555 157.890 8.725 ;
        RECT 157.720 8.195 157.890 8.365 ;
        RECT 150.690 7.475 150.860 7.645 ;
        RECT 150.690 7.115 150.860 7.285 ;
        RECT 150.690 6.755 150.860 6.925 ;
        RECT 150.690 6.395 150.860 6.565 ;
        RECT 150.690 6.035 150.860 6.205 ;
        RECT 150.690 5.675 150.860 5.845 ;
        RECT 150.690 5.315 150.860 5.485 ;
        RECT 150.690 4.955 150.860 5.125 ;
        RECT 150.690 4.595 150.860 4.765 ;
        RECT 152.700 7.720 152.870 7.890 ;
        RECT 153.125 7.720 153.295 7.890 ;
        RECT 153.485 7.720 153.655 7.890 ;
        RECT 153.845 7.720 154.015 7.890 ;
        RECT 154.205 7.720 154.375 7.890 ;
        RECT 154.565 7.720 154.735 7.890 ;
        RECT 154.925 7.720 155.095 7.890 ;
        RECT 155.285 7.720 155.455 7.890 ;
        RECT 155.710 7.720 155.880 7.890 ;
        RECT 152.700 7.295 152.870 7.465 ;
        RECT 152.700 6.935 152.870 7.105 ;
        RECT 155.710 7.295 155.880 7.465 ;
        RECT 155.710 6.935 155.880 7.105 ;
        RECT 152.700 6.575 152.870 6.745 ;
        RECT 152.700 6.215 152.870 6.385 ;
        RECT 152.700 5.855 152.870 6.025 ;
        RECT 153.845 5.855 154.735 6.745 ;
        RECT 155.710 6.575 155.880 6.745 ;
        RECT 155.710 6.215 155.880 6.385 ;
        RECT 155.710 5.855 155.880 6.025 ;
        RECT 152.700 5.495 152.870 5.665 ;
        RECT 152.700 5.135 152.870 5.305 ;
        RECT 155.710 5.495 155.880 5.665 ;
        RECT 155.710 5.135 155.880 5.305 ;
        RECT 152.700 4.710 152.870 4.880 ;
        RECT 153.125 4.710 153.295 4.880 ;
        RECT 153.485 4.710 153.655 4.880 ;
        RECT 153.845 4.710 154.015 4.880 ;
        RECT 154.205 4.710 154.375 4.880 ;
        RECT 154.565 4.710 154.735 4.880 ;
        RECT 154.925 4.710 155.095 4.880 ;
        RECT 155.285 4.710 155.455 4.880 ;
        RECT 155.710 4.710 155.880 4.880 ;
        RECT 157.720 7.835 157.890 8.005 ;
        RECT 157.720 7.475 157.890 7.645 ;
        RECT 157.720 7.115 157.890 7.285 ;
        RECT 157.720 6.755 157.890 6.925 ;
        RECT 157.720 6.395 157.890 6.565 ;
        RECT 157.720 6.035 157.890 6.205 ;
        RECT 157.720 5.675 157.890 5.845 ;
        RECT 157.720 5.315 157.890 5.485 ;
        RECT 157.720 4.955 157.890 5.125 ;
        RECT 150.690 4.235 150.860 4.405 ;
        RECT 150.690 3.875 150.860 4.045 ;
        RECT 150.690 3.515 150.860 3.685 ;
        RECT 150.690 3.155 150.860 3.325 ;
        RECT 157.720 4.595 157.890 4.765 ;
        RECT 157.720 4.235 157.890 4.405 ;
        RECT 157.720 3.875 157.890 4.045 ;
        RECT 157.720 3.515 157.890 3.685 ;
        RECT 157.720 3.155 157.890 3.325 ;
        RECT 150.690 2.700 150.860 2.870 ;
        RECT 151.145 2.700 151.315 2.870 ;
        RECT 151.505 2.700 151.675 2.870 ;
        RECT 151.865 2.700 152.035 2.870 ;
        RECT 152.225 2.700 152.395 2.870 ;
        RECT 152.585 2.700 152.755 2.870 ;
        RECT 152.945 2.700 153.115 2.870 ;
        RECT 153.305 2.700 153.475 2.870 ;
        RECT 153.665 2.700 153.835 2.870 ;
        RECT 154.025 2.700 154.195 2.870 ;
        RECT 154.385 2.700 154.555 2.870 ;
        RECT 154.745 2.700 154.915 2.870 ;
        RECT 155.105 2.700 155.275 2.870 ;
        RECT 155.465 2.700 155.635 2.870 ;
        RECT 155.825 2.700 155.995 2.870 ;
        RECT 156.185 2.700 156.355 2.870 ;
        RECT 156.545 2.700 156.715 2.870 ;
        RECT 156.905 2.700 157.075 2.870 ;
        RECT 157.265 2.700 157.435 2.870 ;
        RECT 157.720 2.700 157.890 2.870 ;
      LAYER met1 ;
        RECT 150.630 9.670 157.950 9.960 ;
        RECT 150.630 2.930 150.920 9.670 ;
        RECT 152.640 7.660 155.940 7.950 ;
        RECT 152.640 4.940 152.930 7.660 ;
        RECT 153.785 5.795 154.795 6.805 ;
        RECT 155.650 4.940 155.940 7.660 ;
        RECT 152.640 4.650 155.940 4.940 ;
        RECT 157.660 2.930 157.950 9.670 ;
        RECT 150.630 2.640 157.950 2.930 ;
  END
END tt_um_example
END LIBRARY

